`include "clk_ibuf.v"
`include "iodelay_ctrl.v"
`include "infrastructure.v"
